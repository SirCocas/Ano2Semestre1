---------------------------------------------------------------------------
-- University of Aveiro - DETI
-- "Computer Architecture I" course (Practical classes)
-- 
-- MIPS multi-cycle datapath
---------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library work;
use work.DisplayUnit_pkg.all;

entity MIPS_MultiCycle is
	port(	clk 			: in std_logic;
			reset			: in std_logic;
			cpu_rd		: out std_logic;
			cpu_wr		: out std_logic;
			cpu_addrBus	: out std_logic_vector(31 downto 0);
			cpu_dataBus	: inout std_logic_vector(31 downto 0)
		);
end MIPS_MultiCycle;

architecture Struct of MIPS_MultiCycle is
-- Signals related to the instruction code
	signal si_instr : std_logic_vector(31 downto 0);
	signal si_opcode, si_funct : std_logic_vector(5 downto 0);
	signal si_rs, si_rt, si_rd, si_writeReg, s_muxM2, s_mux1: std_logic_vector(4 downto 0);
	signal si_imm : std_logic_vector(15 downto 0);
	signal si_jAddr : std_logic_vector(25 downto 0);
	signal si_offset32, si_left2, s_muxM3 : std_logic_vector(31 downto 0);
	
-- Other signals
	signal s_zero : std_logic;
	signal s_pc : std_logic_vector(31 downto 0);
	signal s_aluOper : std_logic_vector(2 downto 0);

-- Data signals
	signal sd_readData1, sd_readData2 : std_logic_vector(31 downto 0);
	signal sd_regA, sd_regB : std_logic_vector(31 downto 0);
	signal sd_aluA, sd_aluB : std_logic_vector(31 downto 0);
	signal sd_aluRes : std_logic_vector(31 downto 0);
	signal sd_aluOut : std_logic_vector(31 downto 0);
	signal sd_data : std_logic_vector(31 downto 0);
	signal sd_writeData : std_logic_vector(31 downto 0);
	
-- Control signals (generated by the control unit)
	signal sc_IorD, sc_RegDst, sc_MemToReg : std_logic;
	signal sc_AluSel_a : std_logic;
	signal sc_AluSel_b, sc_AluOp : std_logic_vector(1 downto 0);	
	signal sc_RegWrite, sc_IrWrite  : std_logic;
	signal sc_PCWrite, sc_PCWriteCond : std_logic;
	signal sc_PCSource : std_logic_vector(1 downto 0);	
	
begin

-- PC update
pcupd:	entity work.PCupdate(Behavioral)	
			---todo not sure if this is right
			port map(clk			=> clk,
						reset			=> reset,
						zero			=> s_zero,
						PCSource		=> sc_PCSource, 
						PCWrite		=> sc_PCWrite,
						PCWriteCond	=> sc_PCWriteCond,
						PC4			=> s_pc,
						BTA			=> sd_aluOut,
						jAddr			=> si_jAddr,
						pc				=> s_pc);

-- MUX M1 (address multiplexer)
mux_m1:	entity work.MUX21_N(Behavioral)
			generic map(N => 32)
			port map(In0	=> s_pc,
						In1	=> sd_aluOut,
						Sel	=> sc_IorD,
						MuxOut=> cpu_addrBus);	-- CPU Address Bus		
					
-- Instruction Register
instReg:	entity work.Register_N(Behavioral)
			port map(clk		=> clk,
						enable	=> sc_IrWrite,
						valIn		=> cpu_dataBus,
						valOut	=> si_instr);

-- Data Register
dataReg:	entity work.Register_N(Behavioral)
			port map(clk		=> clk,
						enable	=> '1',
						valIn		=> cpu_dataBus,	-- CPU Data Bus
						valOut	=> sd_data);
						
-- Splitter
spliter:	entity work.InstSplitter(Behavioral)
			port map(instruction	=> si_instr,
						opcode		=> si_opcode,
						rs				=> si_rs,
						rt				=> si_rt,
						rd				=> si_rd,
						funct			=> si_funct,
						imm			=> si_imm,
						jAddr			=> si_jAddr);

-- MUX M2 (Destination register multiplexer)
mux_m2:	entity work.MUX21_N(Behavioral)
			generic map(N => 5)
			port map(In0	=> si_rt,
						In1	=> si_rd,
						Sel	=> sc_RegDst,
						MuxOut=> s_muxM2);		

-- MUX M3 (Register write data multiplexer)
mux_m3:	entity work.MUX21_N(Behavioral)
			generic map(N => 	32)
			port map(In0	=> sd_aluOut,
						In1	=> sd_data,
						Sel	=> sc_MemToReg,
						MuxOut=> s_muxM3);		
						
-- Register File
regfile:	entity work.RegFile(Structural)
			port map(clk			=> clk,
						writeEnable	=> sc_RegWrite,
						writeReg		=> s_muxM2,
						writeData	=> s_muxM3,
						readReg1		=> si_rs,
						readReg2		=> si_rt,
						readData1	=> sd_readData1,
						readData2	=> sd_readData2);

-- A Register
regA:	entity work.Register_N(Behavioral)
			port map(clk		=> clk,
						enable	=> '1',
						valIn		=> sd_readData1,
						valOut	=> sd_regA);

-- B Register
regB:	entity work.Register_N(Behavioral)
			port map(clk		=> clk,
						enable	=> '1',
						valIn		=> sd_readData2,
						valOut	=> sd_regB);

-- MUX M4 (ALU operand A multiplexer)
mux_m4:	entity work.MUX21_N(Behavioral)
			generic map(N => 32)
			port map(In0	=> s_pc,
						In1	=> sd_regA,
						Sel	=> sc_AluSel_a,
						MuxOut=> sd_aluA);

-- MUX M5 (ALU operand B multiplexer)
mux_m5:	entity work.MUX41_N(Behavioral)
			generic map(N => 32)
			port map(In0	=> sd_regB,
						In1	=> X"00000004",
						In2 	=> si_offset32,
						In3 	=> si_left2,
						Sel	=> sc_AluSel_b,
						MuxOut=> sd_aluB);
						
-- ALU
alu:		entity work.alu32(Behavioral)
			port map(a		=> sd_aluA,
						b  	=> sd_aluB,
						oper	=> s_aluOper,
						res	=> sd_aluRes,
						zero	=> s_zero);
						
-- ALU Control		
alucntl:	entity work.ALUControlUnit(Behavioral)
			port map(ALUop		 => sc_AluOp,
						funct		 => si_funct,
						ALUcontrol=> s_aluOper);
						
-- ALUOut Register
regALU:	entity work.Register_N(Behavioral)
			port map(clk		=> clk,
						enable	=> '1',
						valIn		=> sd_aluRes,
						valOut	=> sd_aluOut);
												
-- left shifter
ls2:		entity work.LeftShifter2(Behavioral)
			port map(dataIn	=> si_offset32,
						dataOut	=> si_left2);
						
-- sign extend
signext:	entity work.SignExtend(Behavioral)
			port map(dataIn	=> si_imm,
						dataOut	=> si_offset32);
						
-- Control Unit											
control:	entity work.ControlUnit(Behavioral)
			port map(Clk			=> clk,
						Reset			=> reset,
						OpCode 		=> si_opcode,
						PCWrite		=> sc_PCWrite,
						IRWrite		=> sc_IrWrite,
						IorD			=> sc_IorD,
						PCSource		=> sc_PCSource,
						RegDest		=> sc_RegDst,
						PCWriteCond	=> sc_PCWriteCond,
						MemRead		=> cpu_rd,			-- CPU read signal
						MemWrite		=> cpu_wr,			-- CPU write signal
						MemToReg		=> sc_MemToReg,
						ALUSelA		=> sc_AluSel_a,
						ALUSelB		=> sc_AluSel_b,
						RegWrite		=> sc_RegWrite,
						ALUop 		=> sc_AluOp);

-- Tri-state logic (data bus)
	cpu_dataBus <= sd_regB when cpu_wr = '1' else (others => 'Z');	-- CPU cpu_dataBus
	
-- Connection to DisplayUnit (ALU result, shown as Instruction Memory Data)
	DU_IMdata <= sd_aluRes;
						
end Struct;

