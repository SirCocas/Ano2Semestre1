---------------------------------------------------------------------------
-- University of Aveiro - DETI
-- "Computer Architecture I" course (Practical classes)
-- 
-- MIPS single-cycle datapath
---------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library work;
use work.DisplayUnit_pkg.all;
use work.MIPS_pkg.all;

entity MIPS_SingleCycle is
	port(	CLOCK_50 : in std_logic;
			KEY  		: in std_logic_vector(3 downto 0);
			SW   		: in std_logic_vector(17 downto 0);
			LEDR  	: out std_logic_vector(17 downto 0);
			LEDG  	: out std_logic_vector(8 downto 0);
			HEX0  	: out std_logic_vector(6 downto 0);
			HEX1  	: out std_logic_vector(6 downto 0);
			HEX2  	: out std_logic_vector(6 downto 0);
			HEX3  	: out std_logic_vector(6 downto 0);
			HEX4  	: out std_logic_vector(6 downto 0);
			HEX5  	: out std_logic_vector(6 downto 0);
			HEX6  	: out std_logic_vector(6 downto 0);
			HEX7  	: out std_logic_vector(6 downto 0));
end MIPS_SingleCycle;

architecture Shell of MIPS_SingleCycle is
-- Data signals
	signal sd_readData1 : std_logic_vector(31 downto 0);
	
-- Control signals (generated by the control unit)
	signal sc_RegDst : std_logic;

-- Signals related to the instruction code
	signal si_instr : std_logic_vector(31 downto 0);

-- Other signals
	signal s_clk : std_logic;
	signal s_pc : std_logic_vector(31 downto 0);
-- Auxiliar
	signal s_jumpAddr: std_logic_vector(25 downto 0);
	signal s_extendImm : std_logic_vector(31 downto 0);
	signal s_immediate: std_logic_vector(15 downto 0);
	signal s_instruction: std_logic_vector(31 downto 0);
	signal s_op: std_logic_vector(5 downto 0);
	signal s_rs: std_logic_vector(4 downto 0);
	signal s_rt: std_logic_vector(4 downto 0);
	signal s_rd: std_logic_vector(4 downto 0);
	signal s_shamt: std_logic_vector(4 downto 0);
	signal s_funct: std_logic_vector(5 downto 0);
	
	
begin

-- PC Update
pcupd:	entity work.PCupdate(Behavioral)	
			port map(clk		=> s_clk,  -- ou KEY[0]?
						reset		=> not KEY(1),
						branch	=> '0',
						jump		=> '0',
						zero		=> '0',
						offset32	=> s_extendImm,
						jAddr26	=> s_jumpAddr,
						pc			=> s_pc);

-- Instruction Memory
instmem:	entity work.InstructionMemory(Behavioral)
			generic map(ADDR_BUS_SIZE => ROM_ADDR_SIZE)
			port map(address		=> s_pc( (ROM_ADDR_SIZE +1) downto 2),  --word adresses! ROM-SIZE = 6 --> 2^6 = words --> 2^6*2^2 = bytes
						readData		=> s_instruction);

-- Splitter
spliter:	entity work.InstrSplitter(Behavioral)
			port map(instruction		=> s_instruction,
						opcode	=> s_op,
						rs			=> s_rs,
						rt			=> s_rt,
						rd			=> s_rd,
						shamt		=> s_shamt,
						funct		=> s_funct,
						imm		=> s_immediate,
						jAddr		=> s_jumpAddr);
	
-- Sign Extender
signext:	entity work.SignExtend(Behavioral)
			port map(dataIn	=> s_immediate,
						dataOut	=> s_extendImm);
	
	--DU_RFdata <= s_instruction;
	DU_DMdata <= (others => '0');	
------------------------------------------------------------------------------
-- Support Modules						
------------------------------------------------------------------------------

-- Display Unit
display:	entity work.DisplayUnit(Behavioral)
			generic map(dataPathType => SINGLE_CYCLE_DP,
							IM_ADDR_SIZE => ROM_ADDR_SIZE,
							DM_ADDR_SIZE => RAM_ADDR_SIZE)
			port map(RefClk	=> CLOCK_50,
						InputSel	=> SW(1 downto 0),	
						DispMode	=> SW(17),
						NextAddr	=> KEY(3),
						Dir		=> KEY(2),
						disp0		=> HEX0,
						disp1		=> HEX1,
						disp2		=> HEX2,
						disp3		=> HEX3,
						disp4		=> HEX4,
						disp5		=> HEX5,
						disp6		=> HEX6,
						disp7		=> HEX7);		

-- Debouncer
debncer:	entity work.DebounceUnit(Behavioral)
			generic map(inPolarity	=> '0',
							outPolarity => '1')
			port map(refClk	=> CLOCK_50, 
						dirtyIn	=> KEY(0), 
						pulsedOut=> s_clk);	
	
	
end Shell;
